`timescale 1ns / 1ps

module hazard_detection_unit(
    input wire [2:0] rs1_ID, rs2_ID,    
    input wire [2:0] rd_EX,             
    input wire MemRead_EX,              
    output wire stall                   
    );
    
    assign stall = 0;

endmodule
