`timescale 1ns / 1ps

module fetch789(
input wire clk,
input wire reset,
input wire flush,
input wire stall,
input wire[7:0]branch_target,
input wire jump,
input wire PC_sel,

output reg[15:0]instruction ,
output reg[7:0] PC_out,
output reg valid
);
 reg [7:0] PC;
 reg halt;
 reg [15:0] instruction_memory [0:255];

    initial begin
        $readmemh("instruction.mem", instruction_memory);
    end
always @(posedge clk or posedge reset)
begin
if(reset)begin
PC_out <= 8'b00;
instruction <= 16'b0;
valid <= 1'b0;
halt <= 1'b0;
end

else if(jump)begin
PC<= instruction[11:4];
end

else if(PC_sel)begin
PC<=branch_target;
end 



else if(flush)begin
PC<=branch_target;
end

else if (halt)begin
valid<=1'b0;
end

else if(instruction_memory[PC][15:12]==4'b1111)begin
halt<=1'b1;
end

else
PC<=PC+1;

end










    
endmodule
